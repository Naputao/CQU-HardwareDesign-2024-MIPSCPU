module controller(
    input wire[5:0] opD,functD,
    output reg jump,
    output reg branch,
    output reg [1:0] alusrc,
    output reg [2:0] regfrom, //000:aluout|001:lw|011:mflo|010:mfhi|100:lb|101:lbu|110:lh|111:lhu //00:w|10:b|11:h
    output reg regwrite,
    output reg regdst,
    output reg [3:0] aluControl,
    output reg isUnsignExt,
    output reg hiRegWrite,
    output reg loRegWrite,
    output reg [1:0] saveReg, //00:no|01:w|10:b|11:h
    output reg id_is_break, id_is_syscall, priorControl, id_is_unfinished
    );
    
    always @(*) begin
        case (opD)
            6'b000000: begin
                case (functD)
                    6'b000000: begin  //sll
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b10;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b000010: begin  //srl
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b10;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1001;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b000011: begin  //sra
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b10;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1010;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b000100: begin  //sllv
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b000110: begin  //srlv
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1001;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b000111: begin  //srav
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1010;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b100000: begin  //add
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0010;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b100001: begin  //addu
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0010;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b100010: begin  //sub
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0110;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b100011: begin  //subu
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0110;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b100100: begin  //and
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b100101: begin  //or
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0001;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b101010: begin  //slt
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0111;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b101011: begin  //sltu
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1101;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b100110: begin  //xor
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1011;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b100111: begin  //nor
                        //20231227
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0011;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b010000: begin      //mfhi
                        saveReg <= 2'b00;
                        regfrom <= 3'b010;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b010010: begin      //mflo
                        saveReg <= 2'b00;
                        regfrom <= 3'b011;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b1;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b010001: begin      //mthi
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b1;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b010011: begin      //mtlo
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b1;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b001000: begin      //jr
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b1;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b001001: begin      //jalr
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b1;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b1;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b011010: begin      //div
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0100;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b011011: begin      //divu
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0101;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b011000: begin      //mult
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1110;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b011001: begin      //multu
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b1111;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b001101: begin      //break
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b1;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    6'b001100: begin      //syscall
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b1;
                        id_is_unfinished <= 1'b0;
                        priorControl <= 1'b0;
                    end
                    default: begin
                        saveReg <= 2'b00;
                        regfrom <= 3'b000;
                        alusrc <= 2'b00;
                        regdst <= 1'b0;
                        regwrite <= 1'b0;
                        branch <= 1'b0;
                        jump <= 1'b0;
                        aluControl <= 4'b0000;
                        isUnsignExt <= 1'b0;
                        hiRegWrite <= 1'b0;
                        loRegWrite <= 1'b0;
                        id_is_break <= 1'b0;
                        id_is_syscall <= 1'b0;
                        id_is_unfinished <= 1'b1;
                        priorControl <= 1'b0;
                    end
                endcase
            end
            6'b010000: begin  // eret, mtc0, mfc0
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b00;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0000;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b1;
            end
            6'b100000: begin       //lb
                //20231227
                saveReg <= 2'b00;
                regfrom <= 3'b100;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b100100: begin       //lbu
                saveReg <= 2'b00;
                regfrom <= 3'b101;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b100001: begin       //lh
                saveReg <= 2'b00;
                regfrom <= 3'b110;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b100101: begin       //lhu
                saveReg <= 2'b00;
                regfrom <= 3'b111;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b100011: begin       //lw
                saveReg <= 2'b00;
                regfrom <= 3'b001;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b101000: begin      //sb
                saveReg <= 2'b10; //00:no|01:w|10:b|11:h
                regfrom <= 3'b000; 
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b101001: begin      //sh
                saveReg <= 2'b11; //00:no|01:w|10:b|11:h
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b101011: begin      //sw
                saveReg <= 2'b01; //00:no|01:w|10:b|11:h
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b000100: begin      //beq
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b00;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b1;
                jump <= 1'b0;
                aluControl <= 4'b0110;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b000101: begin      //bne
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b00;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b1;
                jump <= 1'b0;
                aluControl <= 4'b0110;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b000001: begin      //bgez, bgezal, bltz, bltzal
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b00;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b1;
                jump <= 1'b0;
                aluControl <= 4'b0000;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b000111: begin      //bgtz
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b00;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b1;
                jump <= 1'b0;
                aluControl <= 4'b0110;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b000110: begin      //blez
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b00;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b1;
                jump <= 1'b0;
                aluControl <= 4'b0110;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b001000: begin      //addi
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b001001: begin      //addiu
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0010;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b001010: begin      //slti
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0111;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b001011: begin      //sltiu
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b1101;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b000010: begin      //j
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b00;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b0;
                jump <= 1'b1;
                aluControl <= 4'b0000;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b000011: begin      //jal
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b00;
                regdst <= 1'b1;
                regwrite <= 1'b0;
                branch <= 1'b0;
                jump <= 1'b1;
                aluControl <= 4'b0000;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b001100: begin      //andi
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0000;
                isUnsignExt <= 1'b1;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b001101: begin      //ori
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0001;
                isUnsignExt <= 1'b1;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b001110: begin      //xori
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b1011;
                isUnsignExt <= 1'b1;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            6'b001111: begin      //lui
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b01;
                regdst <= 1'b0;
                regwrite <= 1'b1;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b1100;
                isUnsignExt <= 1'b1;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b0;
                priorControl <= 1'b0;
            end
            default: begin
                saveReg <= 2'b00;
                regfrom <= 3'b000;
                alusrc <= 2'b00;
                regdst <= 1'b0;
                regwrite <= 1'b0;
                branch <= 1'b0;
                jump <= 1'b0;
                aluControl <= 4'b0000;
                isUnsignExt <= 1'b0;
                hiRegWrite <= 1'b0;
                loRegWrite <= 1'b0;
                id_is_break <= 1'b0;
                id_is_syscall <= 1'b0;
                id_is_unfinished <= 1'b1;
                priorControl <= 1'b0;
            end
        endcase
    end
endmodule
